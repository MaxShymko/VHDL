

package funcs is
	
	function next_step (goHome : in boolean, ) return ant_arr is
	begin
		if (goHome = true) then
		  
		else
		  
		end if;
	end next_step;


end funcs;
