package types is

	type ant_arr is array (0 to 1) of integer;

end types;
