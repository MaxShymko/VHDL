entity element is
  port(c1,c2,c3,a1,mc2,mc1: in BIT;
    y2,my2,my1: out BIT);
end element;
architecture struct of element is
component
  mult port(a1,b1,mc2,mc1: in BIT;
  mp2,mp1: out BIT);
end component;
component
  add port(c1,c2,c3: in BIT;
  p2,p1: out BIT);
end component;
signal t: BIT;
begin
  circ1: add port map(c1,c2,c3,y2,t);
  circ2: mult port map(a1,t,mc2,mc1,my2,my1);
end struct;